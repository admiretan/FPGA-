module volleyball(
  input   sys_clk,
  input   sys_rst,
  output  [5:0] sel,
  output  [7:0] seg
  );

endmodule
